library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity ROM is
port(
    addr:in std_logic_vector(7 downto 0);
    clk:in std_logic;
    output:out std_logic_vector(7 downto 0));
end ROM;

architecture behaviour of ROM is
type memory is array ( 0 to 255 ) of std_logic_vector( 7 downto 0 ) ;
constant myrom : memory := (
0 => x"B1" ,1 => x"94" ,2 => x"BA" ,3 => x"C8" ,4 => x"0A" ,5 => x"08" ,6 => x"F5" ,7 => x"3B" , 8 => x"36" ,9 => x"6D" ,10 => x"00" ,11 => x"8E" ,12 => x"58" ,13 => x"4A" ,14 => x"5D" ,15 => x"E4" ,
16 => x"85" ,17 => x"04" ,18 => x"FA" ,19 => x"9D" ,20 => x"1B" ,21 => x"B6" ,22 => x"C7" ,23 => x"AC" ,24 => x"25" ,25 => x"2E" ,26 => x"72" ,27 => x"C2" ,28 => x"02" ,29 => x"FD" ,30 => x"CE" ,31 => x"0D" ,
32 => x"5B" ,33 => x"E3" ,34 => x"D6" ,35 => x"12" ,36 => x"17" ,37 => x"B9" ,38 => x"61" ,39 => x"81" ,40 => x"FE" ,41 => x"67" ,42 => x"86" ,43 => x"AD" ,44 => x"71" ,45 => x"6B" ,46 => x"89" ,47 => x"0B" ,
48 => x"5C" ,49 => x"B0" ,50 => x"C0" ,51 => x"FF" ,52 => x"33" ,53 => x"C3" ,54 => x"56" ,55 => x"B8" ,56 => x"35" ,57 => x"C4" ,58 => x"05" ,59 => x"AE" ,60 => x"D8" ,61 => x"E0" ,62 => x"7F" ,63 => x"99" ,
64 => x"E1" ,65 => x"2B" ,66 => x"DC" ,67 => x"1A" ,68 => x"E2" ,69 => x"82" ,70 => x"57" ,71 => x"EC" ,72 => x"70" ,73 => x"3F" ,74 => x"CC" ,75 => x"F0" ,76 => x"95" ,77 => x"EE" ,78 => x"8D" ,79 => x"F1" ,
80 => x"C1" ,81 => x"AB" ,82 => x"76" ,83 => x"38" ,84 => x"9F" ,85 => x"E6" ,86 => x"78" ,87 => x"CA" ,88 => x"F7" ,89 => x"C6" ,90 => x"F8" ,91 => x"60" ,92 => x"D5" ,93 => x"BB" ,94 => x"9C" ,95 => x"4F" ,
96 => x"F3" ,97 => x"3C" ,98 => x"65" ,99 => x"7B" ,100 => x"63" ,101 => x"7C" ,102 => x"30" ,103 => x"6A" ,104 => x"DD" ,105 => x"4E" ,106 => x"A7" ,107 => x"79" ,108 => x"9E" ,109 => x"B2" ,110 => x"3D" ,111 => x"31" ,
112 => x"3E" ,113 => x"98" ,114 => x"B5" ,115 => x"6E" ,116 => x"27" ,117 => x"D3" ,118 => x"BC" ,119 => x"CF" ,120 => x"59" ,121 => x"1E" ,122 => x"18" ,123 => x"1F" ,124 => x"4C" ,125 => x"5A" ,126 => x"B7" ,127 => x"93" ,
128 => x"E9" ,129 => x"DE" ,130 => x"E7" ,131 => x"2C" ,132 => x"8F" ,133 => x"0C" ,134 => x"0F" ,135 => x"A6" ,136 => x"2D" ,137 => x"DB" ,138 => x"49" ,139 => x"F4" ,140 => x"6F" ,141 => x"73" ,142 => x"96" ,143 => x"47" ,
144 => x"06" ,145 => x"07" ,146 => x"53" ,147 => x"16" ,148 => x"ED" ,149 => x"24" ,150 => x"7A" ,151 => x"37" ,152 => x"39" ,153 => x"CB" ,154 => x"A3" ,155 => x"83" ,156 => x"03" ,157 => x"A9" ,158 => x"8B" ,159 => x"F6" ,
160 => x"92" ,161 => x"BD" ,162 => x"9B" ,163 => x"1C" ,164 => x"E5" ,165 => x"D1" ,166 => x"41" ,167 => x"01" ,168 => x"54" ,169 => x"45" ,170 => x"FB" ,171 => x"C9" ,172 => x"5E" ,173 => x"4D" ,174 => x"0E" ,175 => x"F2" ,
176 => x"68" ,177 => x"20" ,178 => x"80" ,179 => x"AA" ,180 => x"22" ,181 => x"7D" ,182 => x"64" ,183 => x"2F" ,184 => x"26" ,185 => x"87" ,186 => x"F9" ,187 => x"34" ,188 => x"90" ,189 => x"40" ,190 => x"55" ,191 => x"11" ,
192 => x"BE" ,193 => x"32" ,194 => x"97" ,195 => x"13" ,196 => x"43" ,197 => x"FC" ,198 => x"9A" ,199 => x"48" ,200 => x"A0" ,201 => x"2A" ,202 => x"88" ,203 => x"5F" ,204 => x"19" ,205 => x"4B" ,206 => x"09" ,207 => x"A1" ,
208 => x"7E" ,209 => x"CD" ,210 => x"A4" ,211 => x"D0" ,212 => x"15" ,213 => x"44" ,214 => x"AF" ,215 => x"8C" ,216 => x"A5" ,217 => x"84" ,218 => x"50" ,219 => x"BF" ,220 => x"66" ,221 => x"D2" ,222 => x"E8" ,223 => x"8A" ,
224 => x"A2" ,225 => x"D7" ,226 => x"46" ,227 => x"52" ,228 => x"42" ,229 => x"A8" ,230 => x"DF" ,231 => x"B3" ,232 => x"69" ,233 => x"74" ,234 => x"C5" ,235 => x"51" ,236 => x"EB" ,237 => x"23" ,238 => x"29" ,239 => x"21" ,
240 => x"D4" ,241 => x"EF" ,242 => x"D9" ,243 => x"B4" ,244 => x"3A" ,245 => x"62" ,246 => x"28" ,247 => x"75" ,248 => x"91" ,249 => x"14" ,250 => x"10" ,251 => x"EA" ,252 => x"77" ,253 => x"6C" ,254 => x"DA" ,255 => x"1D" ) ;
begin
  process(clk)
    begin
      if(clk='1' and clk'event) then
    output <= myrom(to_integer(unsigned(addr(7 downto 0))));
  end if;
  end process;
end behaviour;